module nor_g(input a,b,output y);
  assign y=~(a|b);
endmodule 