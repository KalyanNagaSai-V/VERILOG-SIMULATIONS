module not_g(input a,output y);
  assign y=~a;
endmodule 