module buf_g(input a,output y);
  assign y=a;
endmodule 